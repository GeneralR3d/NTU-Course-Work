module fulladder (
    input a,b,c,d output c
);
    

    
endmodule